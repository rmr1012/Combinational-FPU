module FPU_tb;

	logic			[31:0] a, b;
	logic				op;
	logic			[31:0]	c;
	logic clk;
	logic rst;

	fp_12 uut(
		.clk(clk), .rst(rst),
		.a(a), .b(b),
		.op(op),
		.c(c)
	);


	initial begin
		op = 0; // add		18 + 17 = 35
		a = 32'b0_10000011_00100000000000000000000; //18
		b = 32'b0_10000011_00010000000000000000000; //17

		//      0_10000100_00011000000000000000000 // resut		nothing outputed, c= is never reached
		#50//#2.5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 1; // subtract	18 - 17 = 1
		#50//#2.5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 0; // add		18 + 17 = 35
		a = 32'b0_10000011_00100000000000000000000; //18
		b = 32'b0_10000011_00010000000000000000000; //17
		//      0_10000100_00011000000000000000000 // resut
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);

		op = 0; // add		18 + (-17) = 1
		a = 32'b01000001100100000000000000000000; //18
		b = 32'b11000001100010000000000000000000; //-17
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 0; // add		-18 + 17 = -1
		a = 32'b11000001100100000000000000000000; //-18
		b = 32'b01000001100010000000000000000000; //17
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 0; // add		-1 + (-1) = -2
		a = 32'b10111111100000000000000000000000; //-1
		b = 32'b10111111100000000000000000000000; //-1
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 1; // subtract	18 - 17 = 1
		a = 32'b01000001100100000000000000000000; // 18
		b = 32'b01000001100010000000000000000000; //17
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 1; // subtract	18 - (-17) = 35
		a = 32'b01000001100100000000000000000000; //18
		b = 32'b11000001100010000000000000000000; //-17
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 1; // subtract	-18 - 17 = -35
		a = 32'b11000001100100000000000000000000; //-18
		b = 32'b01000001100010000000000000000000; //17
		#50//#5
		$display("a:%h  b:%h  c:%h  with op: %h",a,b,c,op);
		op = 1; // subtract	-18 - (-17) = -1
		a = 32'b11000001100100000000000000000000; //-18
		b = 32'b11000001100010000000000000000000; //-17
	end

endmodule
